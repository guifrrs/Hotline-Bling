library ieee;
use ieee.std_logic_1164.all;

entity ROM1 is
  port ( address : in std_logic_vector(4 downto 0);
         data : out std_logic_vector(19 downto 0) );
end entity ROM1;

architecture behavioral of ROM1 is
  type mem is array ( 0 to 2**4 - 1) of std_logic_vector(19 downto 0);
  constant my_Rom : mem := (
    0  => "00000000000000000000", -- Nomes em hexadecimal
    1  => "00000000000000000001",
    2  => "00000000000000000010",
    3  => "00000000000000000011",
    4  => "00000000000000000100",
    5  => "11100000000000000000",
    6  => "11010000000000000000",
    7  => "10110000000000000000",
    8  => "01110000000000000000",
    9  => "11000000000000000000",
    10 => "10010000000000000000",
    11 => "00110000000000000000",
    12 => "10100000000000000000",
    13 => "01010000000000000000",
    14 => "10110010000000000000",
    15 => "11110010000000000000",
begin
   process (address)
   begin
     case address is
       when "00000" => data <= my_rom(0);
       when "00001" => data <= my_rom(1);
       when "00010" => data <= my_rom(2);
       when "00011" => data <= my_rom(3);
       when "00100" => data <= my_rom(4);
       when "00101" => data <= my_rom(5);
       when "00110" => data <= my_rom(6);
       when "00111" => data <= my_rom(7);
       when "01000" => data <= my_rom(8);
       when "01001" => data <= my_rom(9);
       when "01010" => data <= my_rom(10);
       when "01011" => data <= my_rom(11);
       when "01100" => data <= my_rom(12);
       when "01101" => data <= my_rom(13);
       when "01110" => data <= my_rom(14);
       when "01111" => data <= my_rom(15);
       when others => data <= "00000000000000000000"; -- Não mostrar nada
     end case;
  end process;
end architecture behavioral;
